* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                          *
*                                                       *
* Cell Name  : gfet                                     *
* Netlisted  : Fri Aug 23 15:05:31 2013                 *
* PVS Version: 12.1.1-p076 Wed May  1 11:22:57 PDT 2013 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 L(ind_0n4) IND_SEL IND_1(PLUS) IND_1(MINUS)
*.DEVTMPLT 1 L(ind_1n5) IND_SEL IND_2(PLUS) IND_2(MINUS)
*.DEVTMPLT 2 L(ind_2n0) IND_SEL IND_3(PLUS) IND_3(MINUS)
*.DEVTMPLT 3 L(ind_2n8) IND_SEL IND_4(PLUS) IND_4(MINUS)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L PLUS MINUS
.ends L

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: gfet                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt gfet
** N=3 EP=0 FDC=1
M0 3 1 2 gfet W=2e-06 L=1e-06 $X=6000 $Y=4000
.ends gfet
