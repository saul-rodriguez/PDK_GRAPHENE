* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                          *
*                                                       *
* Cell Name  : series_cap                               *
* Netlisted  : Fri Aug 23 12:10:33 2013                 *
* PVS Version: 12.1.1-p076 Wed May  1 11:22:57 PDT 2013 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 L(ind_0n4) IND_SEL IND_1(PLUS) IND_1(MINUS)
*.DEVTMPLT 1 L(ind_1n5) IND_SEL IND_2(PLUS) IND_2(MINUS)
*.DEVTMPLT 2 L(ind_2n0) IND_SEL IND_3(PLUS) IND_3(MINUS)
*.DEVTMPLT 3 L(ind_2n8) IND_SEL IND_4(PLUS) IND_4(MINUS)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L PLUS MINUS
.ends L

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: series_cap                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt series_cap IN OUT
** N=3 EP=2 FDC=2
C0 2 OUT 3.22286e-13 L=1e-05 Er=9.1 TOX=2.5e-08 W=1e-05 $[mim_cap] $X=16400 $Y=34600
C1 IN 2 3.22286e-13 L=1e-05 Er=9.1 TOX=2.5e-08 W=1e-05 $[mim_cap] $X=49800 $Y=34600
.ends series_cap
