* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                          *
*                                                       *
* Cell Name  : test_graph_res_series                    *
* Netlisted  : Fri Aug 23 13:30:14 2013                 *
* PVS Version: 12.1.1-p076 Wed May  1 11:22:57 PDT 2013 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 L(ind_0n4) IND_SEL IND_1(PLUS) IND_1(MINUS)
*.DEVTMPLT 1 L(ind_1n5) IND_SEL IND_2(PLUS) IND_2(MINUS)
*.DEVTMPLT 2 L(ind_2n0) IND_SEL IND_3(PLUS) IND_3(MINUS)
*.DEVTMPLT 3 L(ind_2n8) IND_SEL RES_TER(PLUS) RES_TER(MINUS)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L PLUS MINUS
.ends L

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: test_graph_res_series                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt test_graph_res_series
** N=2 EP=0 FDC=2
X0 1 1 L L=2.8e-09 $[ind_2n8] $X=-9000 $Y=0 $dt=3
X1 1 1 L L=2.8e-09 $[ind_2n8] $X=100000 $Y=0 $dt=3
.ends test_graph_res_series
